////////////////////////////////////////
// DUT /////////////////////////////////
//                                    //
// Go out and do something wonderful. //
//                                    //
////////////////////////////////////////

module dut(
    input logic clk,
    input logic rst
);

////////////////////////////////////////
// Nets ////////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// Logic ///////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// SVAs ////////////////////////////////
////////////////////////////////////////

endmodule
