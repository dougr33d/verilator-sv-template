module top(
    input logic ck,
    input logic rst
);

////////////////////////////////////////
// Nets ////////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// Timeout /////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// DUT /////////////////////////////////
////////////////////////////////////////

dut dut (
    .ck,
    .rst
);

endmodule
