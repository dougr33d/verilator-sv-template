module top(
    input logic clk,
    input logic rst
);

////////////////////////////////////////
// Nets ////////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// Timeout /////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// DUT /////////////////////////////////
////////////////////////////////////////

dut dut (
    .clk,
    .rst
);

endmodule
