`ifndef TOP_SV
`define TOP_SV

module top(
    input logic ck,
    input logic rst
);

////////////////////////////////////////
// Nets ////////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// Timeout /////////////////////////////
////////////////////////////////////////

////////////////////////////////////////
// DUT /////////////////////////////////
////////////////////////////////////////

dut dut (
    .ck,
    .rst
);

endmodule

`endif // TOP_SV
